
library libraryCommon;
use     libraryCommon.P2.all;

entity B1 is

end entity;

architecture rtl of B1 is

begin

end architecture;

