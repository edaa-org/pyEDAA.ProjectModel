
library libraryCommon;
use     libraryCommon.P2.all;

entity A2 is

end entity;

architecture rtl of A2 is

begin
  a : entity work.A1
    port (

    );
end architecture;
