library IEEE;
use     IEEE.std_logic_1164.all;

library libCommon;
use     libCommon.P1.all;

entity A1 is
	port (
		signal Clock : in std_logic
	);
end entity;

architecture rtl of A1 is

begin

end architecture;
