
use work.P1.all;

package P2 is

end package;

package body P2 is

end package body;
