
library libraryCommon;
use     libraryCommon.P1.all;

entity A1 is

end entity;

architecture rtl of A1 is

begin

end architecture;

