
package P1 is

end package;

package body P1 is

end package body;
